`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/07/2018 10:10:33 PM
// Design Name: 
// Module Name: Datapath
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Datapath #(
    parameter PC_W = 9, // Program Counter
    parameter INS_W = 32, // Instruction Width
    parameter RF_ADDRESS = 5, // Register File Address
    parameter DATA_W = 32, // Data WriteData
    parameter DM_ADDRESS = 9, // Data Memory Address
    parameter ALU_CC_W = 4 // ALU Control Code Width
    )(
    input logic clk , reset , // global clock
                              // reset , sets the PC to zero
    RegWrite, MemtoReg,       // Register file writing enable   // Memory or ALU MUX
    ALUsrc2, MemWrite,        // Register file or Immediate MUX // Memory Writing Enable
    MemRead, Branch,          // Memory Reading Enable          // Branch
    ALUsrc1, Jump,            // Register file 1 or PC Mux      // Jump
    input logic [ ALU_CC_W -1:0] ALU_CC, // ALU Control Code ( input of the ALU )
    output logic [6:0] opcode,
    output logic [6:0] Funct7,
    output logic [2:0] Funct3,
    output logic [DATA_W-1:0] WB_Data //ALU_Result
    );

logic [PC_W-1:0] PC, PCPlus4;
logic [PC_W-1:0] PCPlusImm, BranchAddr, Next_PC;
logic [INS_W-1:0] Instr;
logic [DATA_W-1:0] Result;
logic [DATA_W-1:0] Reg1, Reg2;
logic [DATA_W-1:0] ReadData;
logic [DATA_W-1:0] SrcA, SrcB, ALUResult, JumpMuxRes;
logic [DATA_W-1:0] ExtImm;

logic PCSrc; //0: PC+4, 1: Branch address.
logic extendBits;

// next PC
    adder #(9) pcadd (PC, 9'b100, PCPlus4);
    flopr #(9) pcreg (clk, reset, Next_PC, PC);

// branch
    adder #(9) pcaddimm (PC, ExtImm[PC_W-1:0], PCPlusImm);
    mux2 #(9) pcmux (PCPlus4, BranchAddr, (Branch & ~ALUResult[0]), Next_PC); // chooses between pcplus4 and branchaddress  
    mux2 #(9) branchmux (PCPlusImm, ALUResult[PC_W-1:0], Jump, BranchAddr);  // chooses between pcplusimm and aluresult for branchaddr

 //Instruction memory
    instructionmemory instr_mem (PC, Instr);
    
    assign opcode = Instr[6:0];
    assign Funct7 = Instr[31:25];
    assign Funct3 = Instr[14:12];
      
// //Register File
    RegFile rf (clk, reset, RegWrite, Instr[11:7], Instr[19:15], Instr[24:20],
            Result, Reg1, Reg2);
      
    mux2 #(32) resmux (JumpMuxRes, ReadData, MemtoReg, Result);
    mux2 #(32) jumpmux (ALUResult, {23'b0, PCPlus4}, Jump, JumpMuxRes); // stores pc+4 in rd if jump
           
//// sign extend
    imm_Gen Ext_Imm (Instr, ExtImm);

//// ALU
    mux2 #(32) srcamux (Reg1, {23'b0, PC}, ALUsrc1, SrcA);
    mux2 #(32) srcbmux (Reg2, ExtImm, ALUsrc2, SrcB);
    alu alu_module (SrcA, SrcB, ALU_CC, ALUResult);
 
    assign WB_Data = Result;
    
////// Data memory 
	datamemory data_mem (clk, MemRead, MemWrite, Funct3, ALUResult[DM_ADDRESS-1:0], Reg2, ReadData);
     
endmodule